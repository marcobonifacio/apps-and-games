module main

fn main() {
	for val in 0 .. 4 {
		println(val)
	}
}