module main

fn main() {
	mut count := 1
	for {
		println('Hi $count times')
		count += 1
	}
}