module main

fn main() {
	fruits := ['apple', 'banana', 'coconut']
	for idx, ele in fruits {
		println('idx: $idx \t fruit: $ele')
	}
}