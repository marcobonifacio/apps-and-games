module main

fn main() {
	greet := fn (name string) {
		println('Hello, $name')
	}
	greet('Pavan')
	greet('Sahithi')
}